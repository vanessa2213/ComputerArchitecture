package moore_fsm_pkg;

parameter N =  4 ;

typedef enum logic [3:0]{S0, S1, S2, S3, S4, S5, S6, S7, S8, S9}state_d;

endpackage

